library verilog;
use verilog.vl_types.all;
entity read_func is
end read_func;
