library verilog;
use verilog.vl_types.all;
entity all_tb is
end all_tb;
