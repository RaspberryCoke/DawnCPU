library verilog;
use verilog.vl_types.all;
entity read_instr2 is
end read_instr2;
