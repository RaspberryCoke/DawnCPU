library verilog;
use verilog.vl_types.all;
entity fetch_tb is
end fetch_tb;
