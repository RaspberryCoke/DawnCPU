library verilog;
use verilog.vl_types.all;
entity top_single_module is
end top_single_module;
