library verilog;
use verilog.vl_types.all;
entity writeback is
end writeback;
