module writeback(

);

endmodule