library verilog;
use verilog.vl_types.all;
entity read_instr is
end read_instr;
