library verilog;
use verilog.vl_types.all;
entity pc_update_module is
end pc_update_module;
