library verilog;
use verilog.vl_types.all;
entity read2 is
end read2;
