library verilog;
use verilog.vl_types.all;
entity execute_tb is
end execute_tb;
